module setAssociative
(
	input [2:0]  read_address,

	input        set_0_line_0_valid,
	input        set_0_line_0_tag,
	input [15:0] set_0_line_0_block,

	input        set_0_line_1_valid,
	input        set_0_line_1_tag,
	input [15:0] set_0_line_1_block,

	input        set_1_line_0_valid,
	input        set_1_line_0_tag,
	input [15:0] set_1_line_0_block,

	input        set_1_line_1_valid,
	input        set_1_line_1_tag,
	input [15:0] set_1_line_1_block,

	output       read_hit,
	output [7:0] read_byte
);

wire not_read_address_0;

wire set_0_select;
wire set_1_select;

wire set_0_line_0_valid_select;
wire set_0_line_1_valid_select;

wire set_0_line_0_match;
wire set_0_line_1_match;

wire set_0_line_0_valid_select_match;
wire set_0_line_1_valid_select_match;

wire set_0_line_0_valid_match;
wire set_0_line_1_valid_match;
wire set_0_valid_match;

wire set_1_line_0_valid_select;
wire set_1_line_1_valid_select;

wire set_1_line_0_match;
wire set_1_line_1_match;

wire set_1_line_0_valid_select_match;
wire set_1_line_1_valid_select_match;

wire set_1_line_0_valid_match;
wire set_1_line_1_valid_match;
wire set_1_valid_match;

wire set_0_line_0_block_15;
wire set_0_line_0_block_14;
wire set_0_line_0_block_13;
wire set_0_line_0_block_12;
wire set_0_line_0_block_11;
wire set_0_line_0_block_10;
wire set_0_line_0_block_09;
wire set_0_line_0_block_08;
wire set_0_line_0_block_07;
wire set_0_line_0_block_06;
wire set_0_line_0_block_05;
wire set_0_line_0_block_04;
wire set_0_line_0_block_03;
wire set_0_line_0_block_02;
wire set_0_line_0_block_01;
wire set_0_line_0_block_00;

wire set_0_line_0_block_15_match;
wire set_0_line_0_block_14_match;
wire set_0_line_0_block_13_match;
wire set_0_line_0_block_12_match;
wire set_0_line_0_block_11_match;
wire set_0_line_0_block_10_match;
wire set_0_line_0_block_09_match;
wire set_0_line_0_block_08_match;
wire set_0_line_0_block_07_match;
wire set_0_line_0_block_06_match;
wire set_0_line_0_block_05_match;
wire set_0_line_0_block_04_match;
wire set_0_line_0_block_03_match;
wire set_0_line_0_block_02_match;
wire set_0_line_0_block_01_match;
wire set_0_line_0_block_00_match;

wire set_0_line_0_block_15_or_block_07;
wire set_0_line_0_block_14_or_block_06;
wire set_0_line_0_block_13_or_block_05;
wire set_0_line_0_block_12_or_block_04;
wire set_0_line_0_block_11_or_block_03;
wire set_0_line_0_block_10_or_block_02;
wire set_0_line_0_block_09_or_block_01;
wire set_0_line_0_block_08_or_block_00;

wire set_0_line_1_block_15;
wire set_0_line_1_block_14;
wire set_0_line_1_block_13;
wire set_0_line_1_block_12;
wire set_0_line_1_block_11;
wire set_0_line_1_block_10;
wire set_0_line_1_block_09;
wire set_0_line_1_block_08;
wire set_0_line_1_block_07;
wire set_0_line_1_block_06;
wire set_0_line_1_block_05;
wire set_0_line_1_block_04;
wire set_0_line_1_block_03;
wire set_0_line_1_block_02;
wire set_0_line_1_block_01;
wire set_0_line_1_block_00;

wire set_0_line_1_block_15_match;
wire set_0_line_1_block_14_match;
wire set_0_line_1_block_13_match;
wire set_0_line_1_block_12_match;
wire set_0_line_1_block_11_match;
wire set_0_line_1_block_10_match;
wire set_0_line_1_block_09_match;
wire set_0_line_1_block_08_match;
wire set_0_line_1_block_07_match;
wire set_0_line_1_block_06_match;
wire set_0_line_1_block_05_match;
wire set_0_line_1_block_04_match;
wire set_0_line_1_block_03_match;
wire set_0_line_1_block_02_match;
wire set_0_line_1_block_01_match;
wire set_0_line_1_block_00_match;

wire set_0_line_1_block_15_or_block_07;
wire set_0_line_1_block_14_or_block_06;
wire set_0_line_1_block_13_or_block_05;
wire set_0_line_1_block_12_or_block_04;
wire set_0_line_1_block_11_or_block_03;
wire set_0_line_1_block_10_or_block_02;
wire set_0_line_1_block_09_or_block_01;
wire set_0_line_1_block_08_or_block_00;

wire set_0_block_07;
wire set_0_block_06;
wire set_0_block_05;
wire set_0_block_04;
wire set_0_block_03;
wire set_0_block_02;
wire set_0_block_01;
wire set_0_block_00;

wire set_1_line_0_block_15;
wire set_1_line_0_block_14;
wire set_1_line_0_block_13;
wire set_1_line_0_block_12;
wire set_1_line_0_block_11;
wire set_1_line_0_block_10;
wire set_1_line_0_block_09;
wire set_1_line_0_block_08;
wire set_1_line_0_block_07;
wire set_1_line_0_block_06;
wire set_1_line_0_block_05;
wire set_1_line_0_block_04;
wire set_1_line_0_block_03;
wire set_1_line_0_block_02;
wire set_1_line_0_block_01;
wire set_1_line_0_block_00;

wire set_1_line_0_block_15_match;
wire set_1_line_0_block_14_match;
wire set_1_line_0_block_13_match;
wire set_1_line_0_block_12_match;
wire set_1_line_0_block_11_match;
wire set_1_line_0_block_10_match;
wire set_1_line_0_block_09_match;
wire set_1_line_0_block_08_match;
wire set_1_line_0_block_07_match;
wire set_1_line_0_block_06_match;
wire set_1_line_0_block_05_match;
wire set_1_line_0_block_04_match;
wire set_1_line_0_block_03_match;
wire set_1_line_0_block_02_match;
wire set_1_line_0_block_01_match;
wire set_1_line_0_block_00_match;

wire set_1_line_0_block_15_or_block_07;
wire set_1_line_0_block_14_or_block_06;
wire set_1_line_0_block_13_or_block_05;
wire set_1_line_0_block_12_or_block_04;
wire set_1_line_0_block_11_or_block_03;
wire set_1_line_0_block_10_or_block_02;
wire set_1_line_0_block_09_or_block_01;
wire set_1_line_0_block_08_or_block_00;

wire set_1_line_1_block_15;
wire set_1_line_1_block_14;
wire set_1_line_1_block_13;
wire set_1_line_1_block_12;
wire set_1_line_1_block_11;
wire set_1_line_1_block_10;
wire set_1_line_1_block_09;
wire set_1_line_1_block_08;
wire set_1_line_1_block_07;
wire set_1_line_1_block_06;
wire set_1_line_1_block_05;
wire set_1_line_1_block_04;
wire set_1_line_1_block_03;
wire set_1_line_1_block_02;
wire set_1_line_1_block_01;
wire set_1_line_1_block_00;

wire set_1_line_1_block_15_match;
wire set_1_line_1_block_14_match;
wire set_1_line_1_block_13_match;
wire set_1_line_1_block_12_match;
wire set_1_line_1_block_11_match;
wire set_1_line_1_block_10_match;
wire set_1_line_1_block_09_match;
wire set_1_line_1_block_08_match;
wire set_1_line_1_block_07_match;
wire set_1_line_1_block_06_match;
wire set_1_line_1_block_05_match;
wire set_1_line_1_block_04_match;
wire set_1_line_1_block_03_match;
wire set_1_line_1_block_02_match;
wire set_1_line_1_block_01_match;
wire set_1_line_1_block_00_match;

wire set_1_line_1_block_15_or_block_07;
wire set_1_line_1_block_14_or_block_06;
wire set_1_line_1_block_13_or_block_05;
wire set_1_line_1_block_12_or_block_04;
wire set_1_line_1_block_11_or_block_03;
wire set_1_line_1_block_10_or_block_02;
wire set_1_line_1_block_09_or_block_01;
wire set_1_line_1_block_08_or_block_00;

wire set_1_block_07;
wire set_1_block_06;
wire set_1_block_05;
wire set_1_block_04;
wire set_1_block_03;
wire set_1_block_02;
wire set_1_block_01;
wire set_1_block_00;

assign not_read_address_0 = ~ read_address[0];

assign set_0_select = ~ read_address[1];
assign set_1_select =   read_address[1];

assign set_0_line_0_valid_select = set_0_select & set_0_line_0_valid;
assign set_0_line_1_valid_select = set_0_select & set_0_line_1_valid;

assign set_0_line_0_match = read_address[2] ~^ set_0_line_0_tag;
assign set_0_line_1_match = read_address[2] ~^ set_0_line_1_tag;

assign set_0_line_0_valid_select_match = set_0_line_0_valid_select & set_0_line_0_match;
assign set_0_line_1_valid_select_match = set_0_line_1_valid_select & set_0_line_1_match;

assign set_0_line_0_valid_match = set_0_select & set_0_line_0_match;
assign set_0_line_1_valid_match = set_0_select & set_0_line_1_match;

assign set_0_valid_match = set_0_line_0_valid_select_match | set_0_line_1_valid_select_match;

assign set_1_line_0_valid_select = set_1_select & set_1_line_0_valid;
assign set_1_line_1_valid_select = set_1_select & set_1_line_1_valid;

assign set_1_line_0_match = read_address[2] ~^ set_1_line_0_tag;
assign set_1_line_1_match = read_address[2] ~^ set_1_line_1_tag;

assign set_1_line_0_valid_select_match = set_1_line_0_valid_select & set_1_line_0_match;
assign set_1_line_1_valid_select_match = set_1_line_1_valid_select & set_1_line_1_match;

assign set_1_line_0_valid_match = set_1_select & set_1_line_0_match;
assign set_1_line_1_valid_match = set_1_select & set_1_line_1_match;

assign set_1_valid_match = set_1_line_0_valid_select_match | set_1_line_1_valid_select_match;

assign read_hit = set_0_valid_match | set_1_valid_match;

assign set_0_line_0_block_15 = read_address[0] & set_0_line_0_block[15];
assign set_0_line_0_block_14 = read_address[0] & set_0_line_0_block[14];
assign set_0_line_0_block_13 = read_address[0] & set_0_line_0_block[13];
assign set_0_line_0_block_12 = read_address[0] & set_0_line_0_block[12];
assign set_0_line_0_block_11 = read_address[0] & set_0_line_0_block[11];
assign set_0_line_0_block_10 = read_address[0] & set_0_line_0_block[10];
assign set_0_line_0_block_09 = read_address[0] & set_0_line_0_block[9];
assign set_0_line_0_block_08 = read_address[0] & set_0_line_0_block[8];
assign set_0_line_0_block_07 = not_read_address_0 & set_0_line_0_block[7];
assign set_0_line_0_block_06 = not_read_address_0 & set_0_line_0_block[6];
assign set_0_line_0_block_05 = not_read_address_0 & set_0_line_0_block[5];
assign set_0_line_0_block_04 = not_read_address_0 & set_0_line_0_block[4];
assign set_0_line_0_block_03 = not_read_address_0 & set_0_line_0_block[3];
assign set_0_line_0_block_02 = not_read_address_0 & set_0_line_0_block[2];
assign set_0_line_0_block_01 = not_read_address_0 & set_0_line_0_block[1];
assign set_0_line_0_block_00 = not_read_address_0 & set_0_line_0_block[0];

assign set_0_line_0_block_15_match = set_0_line_0_valid_match & set_0_line_0_block_15;
assign set_0_line_0_block_14_match = set_0_line_0_valid_match & set_0_line_0_block_14;
assign set_0_line_0_block_13_match = set_0_line_0_valid_match & set_0_line_0_block_13;
assign set_0_line_0_block_12_match = set_0_line_0_valid_match & set_0_line_0_block_12;
assign set_0_line_0_block_11_match = set_0_line_0_valid_match & set_0_line_0_block_11;
assign set_0_line_0_block_10_match = set_0_line_0_valid_match & set_0_line_0_block_10;
assign set_0_line_0_block_09_match = set_0_line_0_valid_match & set_0_line_0_block_09;
assign set_0_line_0_block_08_match = set_0_line_0_valid_match & set_0_line_0_block_08;
assign set_0_line_0_block_07_match = set_0_line_0_valid_match & set_0_line_0_block_07;
assign set_0_line_0_block_06_match = set_0_line_0_valid_match & set_0_line_0_block_06;
assign set_0_line_0_block_05_match = set_0_line_0_valid_match & set_0_line_0_block_05;
assign set_0_line_0_block_04_match = set_0_line_0_valid_match & set_0_line_0_block_04;
assign set_0_line_0_block_03_match = set_0_line_0_valid_match & set_0_line_0_block_03;
assign set_0_line_0_block_02_match = set_0_line_0_valid_match & set_0_line_0_block_02;
assign set_0_line_0_block_01_match = set_0_line_0_valid_match & set_0_line_0_block_01;
assign set_0_line_0_block_00_match = set_0_line_0_valid_match & set_0_line_0_block_00;

assign set_0_line_0_block_15_or_block_07 = set_0_line_0_block_15_match | set_0_line_0_block_07_match;
assign set_0_line_0_block_14_or_block_06 = set_0_line_0_block_14_match | set_0_line_0_block_06_match;
assign set_0_line_0_block_13_or_block_05 = set_0_line_0_block_13_match | set_0_line_0_block_05_match;
assign set_0_line_0_block_12_or_block_04 = set_0_line_0_block_12_match | set_0_line_0_block_04_match;
assign set_0_line_0_block_11_or_block_03 = set_0_line_0_block_11_match | set_0_line_0_block_03_match;
assign set_0_line_0_block_10_or_block_02 = set_0_line_0_block_10_match | set_0_line_0_block_02_match;
assign set_0_line_0_block_09_or_block_01 = set_0_line_0_block_09_match | set_0_line_0_block_01_match;
assign set_0_line_0_block_08_or_block_00 = set_0_line_0_block_08_match | set_0_line_0_block_00_match;

assign set_0_line_1_block_15 = read_address[0] & set_0_line_1_block[15];
assign set_0_line_1_block_14 = read_address[0] & set_0_line_1_block[14];
assign set_0_line_1_block_13 = read_address[0] & set_0_line_1_block[13];
assign set_0_line_1_block_12 = read_address[0] & set_0_line_1_block[12];
assign set_0_line_1_block_11 = read_address[0] & set_0_line_1_block[11];
assign set_0_line_1_block_10 = read_address[0] & set_0_line_1_block[10];
assign set_0_line_1_block_09 = read_address[0] & set_0_line_1_block[9];
assign set_0_line_1_block_08 = read_address[0] & set_0_line_1_block[8];
assign set_0_line_1_block_07 = not_read_address_0 & set_0_line_1_block[7];
assign set_0_line_1_block_06 = not_read_address_0 & set_0_line_1_block[6];
assign set_0_line_1_block_05 = not_read_address_0 & set_0_line_1_block[5];
assign set_0_line_1_block_04 = not_read_address_0 & set_0_line_1_block[4];
assign set_0_line_1_block_03 = not_read_address_0 & set_0_line_1_block[3];
assign set_0_line_1_block_02 = not_read_address_0 & set_0_line_1_block[2];
assign set_0_line_1_block_01 = not_read_address_0 & set_0_line_1_block[1];
assign set_0_line_1_block_00 = not_read_address_0 & set_0_line_1_block[0];

assign set_0_line_1_block_15_match = set_0_line_1_valid_match & set_0_line_1_block_15;
assign set_0_line_1_block_14_match = set_0_line_1_valid_match & set_0_line_1_block_14;
assign set_0_line_1_block_13_match = set_0_line_1_valid_match & set_0_line_1_block_13;
assign set_0_line_1_block_12_match = set_0_line_1_valid_match & set_0_line_1_block_12;
assign set_0_line_1_block_11_match = set_0_line_1_valid_match & set_0_line_1_block_11;
assign set_0_line_1_block_10_match = set_0_line_1_valid_match & set_0_line_1_block_10;
assign set_0_line_1_block_09_match = set_0_line_1_valid_match & set_0_line_1_block_09;
assign set_0_line_1_block_08_match = set_0_line_1_valid_match & set_0_line_1_block_08;
assign set_0_line_1_block_07_match = set_0_line_1_valid_match & set_0_line_1_block_07;
assign set_0_line_1_block_06_match = set_0_line_1_valid_match & set_0_line_1_block_06;
assign set_0_line_1_block_05_match = set_0_line_1_valid_match & set_0_line_1_block_05;
assign set_0_line_1_block_04_match = set_0_line_1_valid_match & set_0_line_1_block_04;
assign set_0_line_1_block_03_match = set_0_line_1_valid_match & set_0_line_1_block_03;
assign set_0_line_1_block_02_match = set_0_line_1_valid_match & set_0_line_1_block_02;
assign set_0_line_1_block_01_match = set_0_line_1_valid_match & set_0_line_1_block_01;
assign set_0_line_1_block_00_match = set_0_line_1_valid_match & set_0_line_1_block_00;

assign set_0_line_1_block_15_or_block_07 = set_0_line_1_block_15_match | set_0_line_1_block_07_match;
assign set_0_line_1_block_14_or_block_06 = set_0_line_1_block_14_match | set_0_line_1_block_06_match;
assign set_0_line_1_block_13_or_block_05 = set_0_line_1_block_13_match | set_0_line_1_block_05_match;
assign set_0_line_1_block_12_or_block_04 = set_0_line_1_block_12_match | set_0_line_1_block_04_match;
assign set_0_line_1_block_11_or_block_03 = set_0_line_1_block_11_match | set_0_line_1_block_03_match;
assign set_0_line_1_block_10_or_block_02 = set_0_line_1_block_10_match | set_0_line_1_block_02_match;
assign set_0_line_1_block_09_or_block_01 = set_0_line_1_block_09_match | set_0_line_1_block_01_match;
assign set_0_line_1_block_08_or_block_00 = set_0_line_1_block_08_match | set_0_line_1_block_00_match;

assign set_0_block_07 = set_0_line_0_block_15_or_block_07 | set_0_line_1_block_15_or_block_07;
assign set_0_block_06 = set_0_line_0_block_14_or_block_06 | set_0_line_1_block_14_or_block_06;
assign set_0_block_05 = set_0_line_0_block_13_or_block_05 | set_0_line_1_block_13_or_block_05;
assign set_0_block_04 = set_0_line_0_block_12_or_block_04 | set_0_line_1_block_12_or_block_04;
assign set_0_block_03 = set_0_line_0_block_11_or_block_03 | set_0_line_1_block_11_or_block_03;
assign set_0_block_02 = set_0_line_0_block_10_or_block_02 | set_0_line_1_block_10_or_block_02;
assign set_0_block_01 = set_0_line_0_block_09_or_block_01 | set_0_line_1_block_09_or_block_01;
assign set_0_block_00 = set_0_line_0_block_08_or_block_00 | set_0_line_1_block_08_or_block_00;

assign set_1_line_0_block_15 = read_address[0] & set_1_line_0_block[15];
assign set_1_line_0_block_14 = read_address[0] & set_1_line_0_block[14];
assign set_1_line_0_block_13 = read_address[0] & set_1_line_0_block[13];
assign set_1_line_0_block_12 = read_address[0] & set_1_line_0_block[12];
assign set_1_line_0_block_11 = read_address[0] & set_1_line_0_block[11];
assign set_1_line_0_block_10 = read_address[0] & set_1_line_0_block[10];
assign set_1_line_0_block_09 = read_address[0] & set_1_line_0_block[9];
assign set_1_line_0_block_08 = read_address[0] & set_1_line_0_block[8];
assign set_1_line_0_block_07 = not_read_address_0 & set_1_line_0_block[7];
assign set_1_line_0_block_06 = not_read_address_0 & set_1_line_0_block[6];
assign set_1_line_0_block_05 = not_read_address_0 & set_1_line_0_block[5];
assign set_1_line_0_block_04 = not_read_address_0 & set_1_line_0_block[4];
assign set_1_line_0_block_03 = not_read_address_0 & set_1_line_0_block[3];
assign set_1_line_0_block_02 = not_read_address_0 & set_1_line_0_block[2];
assign set_1_line_0_block_01 = not_read_address_0 & set_1_line_0_block[1];
assign set_1_line_0_block_00 = not_read_address_0 & set_1_line_0_block[0];

assign set_1_line_0_block_15_match = set_1_line_0_valid_match & set_1_line_0_block_15;
assign set_1_line_0_block_14_match = set_1_line_0_valid_match & set_1_line_0_block_14;
assign set_1_line_0_block_13_match = set_1_line_0_valid_match & set_1_line_0_block_13;
assign set_1_line_0_block_12_match = set_1_line_0_valid_match & set_1_line_0_block_12;
assign set_1_line_0_block_11_match = set_1_line_0_valid_match & set_1_line_0_block_11;
assign set_1_line_0_block_10_match = set_1_line_0_valid_match & set_1_line_0_block_10;
assign set_1_line_0_block_09_match = set_1_line_0_valid_match & set_1_line_0_block_09;
assign set_1_line_0_block_08_match = set_1_line_0_valid_match & set_1_line_0_block_08;
assign set_1_line_0_block_07_match = set_1_line_0_valid_match & set_1_line_0_block_07;
assign set_1_line_0_block_06_match = set_1_line_0_valid_match & set_1_line_0_block_06;
assign set_1_line_0_block_05_match = set_1_line_0_valid_match & set_1_line_0_block_05;
assign set_1_line_0_block_04_match = set_1_line_0_valid_match & set_1_line_0_block_04;
assign set_1_line_0_block_03_match = set_1_line_0_valid_match & set_1_line_0_block_03;
assign set_1_line_0_block_02_match = set_1_line_0_valid_match & set_1_line_0_block_02;
assign set_1_line_0_block_01_match = set_1_line_0_valid_match & set_1_line_0_block_01;
assign set_1_line_0_block_00_match = set_1_line_0_valid_match & set_1_line_0_block_00;

assign set_1_line_0_block_15_or_block_07 = set_1_line_0_block_15_match | set_1_line_0_block_07_match;
assign set_1_line_0_block_14_or_block_06 = set_1_line_0_block_14_match | set_1_line_0_block_06_match;
assign set_1_line_0_block_13_or_block_05 = set_1_line_0_block_13_match | set_1_line_0_block_05_match;
assign set_1_line_0_block_12_or_block_04 = set_1_line_0_block_12_match | set_1_line_0_block_04_match;
assign set_1_line_0_block_11_or_block_03 = set_1_line_0_block_11_match | set_1_line_0_block_03_match;
assign set_1_line_0_block_10_or_block_02 = set_1_line_0_block_10_match | set_1_line_0_block_02_match;
assign set_1_line_0_block_09_or_block_01 = set_1_line_0_block_09_match | set_1_line_0_block_01_match;
assign set_1_line_0_block_08_or_block_00 = set_1_line_0_block_08_match | set_1_line_0_block_00_match;

assign set_1_line_1_block_15 = read_address[0] & set_1_line_1_block[15];
assign set_1_line_1_block_14 = read_address[0] & set_1_line_1_block[14];
assign set_1_line_1_block_13 = read_address[0] & set_1_line_1_block[13];
assign set_1_line_1_block_12 = read_address[0] & set_1_line_1_block[12];
assign set_1_line_1_block_11 = read_address[0] & set_1_line_1_block[11];
assign set_1_line_1_block_10 = read_address[0] & set_1_line_1_block[10];
assign set_1_line_1_block_09 = read_address[0] & set_1_line_1_block[9];
assign set_1_line_1_block_08 = read_address[0] & set_1_line_1_block[8];
assign set_1_line_1_block_07 = not_read_address_0 & set_1_line_1_block[7];
assign set_1_line_1_block_06 = not_read_address_0 & set_1_line_1_block[6];
assign set_1_line_1_block_05 = not_read_address_0 & set_1_line_1_block[5];
assign set_1_line_1_block_04 = not_read_address_0 & set_1_line_1_block[4];
assign set_1_line_1_block_03 = not_read_address_0 & set_1_line_1_block[3];
assign set_1_line_1_block_02 = not_read_address_0 & set_1_line_1_block[2];
assign set_1_line_1_block_01 = not_read_address_0 & set_1_line_1_block[1];
assign set_1_line_1_block_00 = not_read_address_0 & set_1_line_1_block[0];

assign set_1_line_1_block_15_match = set_1_line_1_valid_match & set_1_line_1_block_15;
assign set_1_line_1_block_14_match = set_1_line_1_valid_match & set_1_line_1_block_14;
assign set_1_line_1_block_13_match = set_1_line_1_valid_match & set_1_line_1_block_13;
assign set_1_line_1_block_12_match = set_1_line_1_valid_match & set_1_line_1_block_12;
assign set_1_line_1_block_11_match = set_1_line_1_valid_match & set_1_line_1_block_11;
assign set_1_line_1_block_10_match = set_1_line_1_valid_match & set_1_line_1_block_10;
assign set_1_line_1_block_09_match = set_1_line_1_valid_match & set_1_line_1_block_09;
assign set_1_line_1_block_08_match = set_1_line_1_valid_match & set_1_line_1_block_08;
assign set_1_line_1_block_07_match = set_1_line_1_valid_match & set_1_line_1_block_07;
assign set_1_line_1_block_06_match = set_1_line_1_valid_match & set_1_line_1_block_06;
assign set_1_line_1_block_05_match = set_1_line_1_valid_match & set_1_line_1_block_05;
assign set_1_line_1_block_04_match = set_1_line_1_valid_match & set_1_line_1_block_04;
assign set_1_line_1_block_03_match = set_1_line_1_valid_match & set_1_line_1_block_03;
assign set_1_line_1_block_02_match = set_1_line_1_valid_match & set_1_line_1_block_02;
assign set_1_line_1_block_01_match = set_1_line_1_valid_match & set_1_line_1_block_01;
assign set_1_line_1_block_00_match = set_1_line_1_valid_match & set_1_line_1_block_00;

assign set_1_line_1_block_15_or_block_07 = set_1_line_1_block_15_match | set_1_line_1_block_07_match;
assign set_1_line_1_block_14_or_block_06 = set_1_line_1_block_14_match | set_1_line_1_block_06_match;
assign set_1_line_1_block_13_or_block_05 = set_1_line_1_block_13_match | set_1_line_1_block_05_match;
assign set_1_line_1_block_12_or_block_04 = set_1_line_1_block_12_match | set_1_line_1_block_04_match;
assign set_1_line_1_block_11_or_block_03 = set_1_line_1_block_11_match | set_1_line_1_block_03_match;
assign set_1_line_1_block_10_or_block_02 = set_1_line_1_block_10_match | set_1_line_1_block_02_match;
assign set_1_line_1_block_09_or_block_01 = set_1_line_1_block_09_match | set_1_line_1_block_01_match;
assign set_1_line_1_block_08_or_block_00 = set_1_line_1_block_08_match | set_1_line_1_block_00_match;

assign set_1_block_07 = set_1_line_0_block_15_or_block_07 | set_1_line_1_block_15_or_block_07;
assign set_1_block_06 = set_1_line_0_block_14_or_block_06 | set_1_line_1_block_14_or_block_06;
assign set_1_block_05 = set_1_line_0_block_13_or_block_05 | set_1_line_1_block_13_or_block_05;
assign set_1_block_04 = set_1_line_0_block_12_or_block_04 | set_1_line_1_block_12_or_block_04;
assign set_1_block_03 = set_1_line_0_block_11_or_block_03 | set_1_line_1_block_11_or_block_03;
assign set_1_block_02 = set_1_line_0_block_10_or_block_02 | set_1_line_1_block_10_or_block_02;
assign set_1_block_01 = set_1_line_0_block_09_or_block_01 | set_1_line_1_block_09_or_block_01;
assign set_1_block_00 = set_1_line_0_block_08_or_block_00 | set_1_line_1_block_08_or_block_00;

assign read_byte[7] = set_0_block_07 | set_1_block_07;
assign read_byte[6] = set_0_block_06 | set_1_block_06;
assign read_byte[5] = set_0_block_05 | set_1_block_05;
assign read_byte[4] = set_0_block_04 | set_1_block_04;
assign read_byte[3] = set_0_block_03 | set_1_block_03;
assign read_byte[2] = set_0_block_02 | set_1_block_02;
assign read_byte[1] = set_0_block_01 | set_1_block_01;
assign read_byte[0] = set_0_block_00 | set_1_block_00;
endmodule
